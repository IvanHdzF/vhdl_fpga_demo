library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity tb_spi_slave_phy is
end entity tb_spi_slave_phy;

architecture sim of tb_spi_slave_phy is

  -- DUT ports
  signal sclk    : std_logic := '0';
  signal cs_n    : std_logic := '1';
  signal mosi    : std_logic := '0';
  signal miso    : std_logic;

  signal rx_byte  : std_logic_vector(7 downto 0);
  signal rx_valid : std_logic;
  signal tx_byte  : std_logic_vector(7 downto 0) := (others => '0');
  signal tx_valid : std_logic := '0';
  signal tx_ready : std_logic;

  constant C_SCLK_PERIOD : time := 20 ns;

begin

  ---------------------------------------------------------------------------
  -- Instantiate DUT
  ---------------------------------------------------------------------------
  dut : entity work.spi_slave_phy
    generic map (
      G_CPOL => '0',
      G_CPHA => '0'
    )
    port map (
      sclk     => sclk,
      cs_n     => cs_n,
      mosi     => mosi,
      miso     => miso,
      rx_byte  => rx_byte,
      rx_valid => rx_valid,
      tx_byte  => tx_byte,
      tx_valid => tx_valid,
      tx_ready => tx_ready
    );

  ---------------------------------------------------------------------------
  -- Generate SCLK
  ---------------------------------------------------------------------------
  sclk_gen : process
  begin
    while true loop
      sclk <= '0';
      wait for C_SCLK_PERIOD/2;
      sclk <= '1';
      wait for C_SCLK_PERIOD/2;
    end loop;
  end process;

  ---------------------------------------------------------------------------
  -- Stimulus process
  ---------------------------------------------------------------------------
  stim : process
    procedure spi_send_byte(constant b : std_logic_vector(7 downto 0)) is
    begin
      -- MSB first, change MOSI on falling, sample on rising (mode 0)
      for i in 7 downto 0 loop
        wait until falling_edge(sclk);
        mosi <= b(i);
        wait until rising_edge(sclk);
      end loop;
    end procedure;

    -- Full-duplex: send one byte on MOSI, capture one byte from MISO
    procedure spi_full_duplex(
      constant mosi_byte : std_logic_vector(7 downto 0);
      variable miso_byte : out std_logic_vector(7 downto 0)
    ) is
    begin
      for i in 7 downto 0 loop
        wait until falling_edge(sclk);
        mosi <= mosi_byte(i);      -- master drives MOSI
        wait until rising_edge(sclk);
        miso_byte(i) := miso;      -- master samples MISO
      end loop;
    end procedure;

    -- local variables
    variable tx_sampled  : std_logic_vector(7 downto 0);
    variable tx_sampled2 : std_logic_vector(7 downto 0);
    variable error_count : integer := 0;

     -- for multi-byte full-duplex test
    type t_byte_arr is array (0 to 3) of std_logic_vector(7 downto 0);
    variable mosi_seq    : t_byte_arr := (x"A1", x"B2", x"C3", x"D4");
    variable miso_seq    : t_byte_arr := (x"11", x"22", x"33", x"44");
    variable mosi_captured : t_byte_arr;
    variable miso_captured : t_byte_arr;

  begin
    -- Initial idle
    cs_n    <= '1';
    mosi    <= '0';
    tx_byte <= (others => '0');
    tx_valid<= '0';
    wait for 5*C_SCLK_PERIOD;

    -------------------------------------------------------------------------
    -- Test 1: RX only, send 0xF0 from master to slave
    -------------------------------------------------------------------------
    report "Test 1: RX path, sending 0xF0" severity note;
    cs_n <= '0';
    spi_send_byte(x"F0");

    -- Wait for full byte
    wait until rx_valid = '1';
    wait until falling_edge(sclk);  -- settle

    if rx_byte /= x"F0" then
      error_count := error_count + 1;
      report "Test 1 FAILED. rx_byte dec=" &
             integer'image(to_integer(unsigned(rx_byte)))
        severity error;
    else
      report "Test 1 PASSED" severity note;
    end if;

    wait until rising_edge(sclk);
    cs_n <= '1';
    wait for C_SCLK_PERIOD;  -- CS high ≥ 1 SCLK
    wait for C_SCLK_PERIOD;

    mosi <= '0';

    -------------------------------------------------------------------------
    -- Test 2: TX path, have slave transmit 0x5A while master clocks
    -------------------------------------------------------------------------
    report "Test 2: TX path, transmitting 0x5A" severity note;
    tx_byte  <= x"5A";
    tx_valid <= '1';  -- DUT will sample when tx_ready='1'

    tx_sampled := (others => '0');

    cs_n <= '0';
    -- Slave updates MISO on falling; master samples on rising
    for i in 7 downto 0 loop
      wait until falling_edge(sclk);
      
      wait until rising_edge(sclk);
      tx_sampled(i) := miso;
      report "MISO bit index " & integer'image(i) &
             " = " & std_logic'image(miso)
        severity note;
    end loop;
    cs_n <= '1';
    tx_valid <= '0';
    wait until falling_edge(sclk);
    wait for C_SCLK_PERIOD;  -- CS high ≥ 1 SCLK
    wait for C_SCLK_PERIOD;

    if tx_sampled /= x"5A" then
      error_count := error_count + 1;
      report "Test 2 FAILED. tx_sampled dec=" &
             integer'image(to_integer(unsigned(tx_sampled)))
        severity error;
    else
      report "Test 2 PASSED" severity note;
    end if;

    -------------------------------------------------------------------------
    -- Test 3: Full-duplex, 1 byte RX + 1 byte TX in same CS
    -------------------------------------------------------------------------
    report "Test 3: Full-duplex, RX 0xA5 while TX 0x3C" severity note;

    tx_byte  <= x"3C";
    tx_valid <= '1';
    tx_sampled := (others => '0');
    cs_n <= '0';

    -- send 0xA5 on MOSI, capture MISO simultaneously
    spi_full_duplex(x"A5", tx_sampled);

    -- Wait for rx_valid and settle
    wait until rx_valid = '1';
    wait until falling_edge(sclk);

    -- end of frame
    cs_n <= '1';
    tx_valid <= '0';

    if rx_byte /= x"A5" then
      error_count := error_count + 1;
      report "Test 3 FAILED RX. rx_byte dec=" &
             integer'image(to_integer(unsigned(rx_byte)))
        severity error;
    elsif tx_sampled /= x"3C" then
      error_count := error_count + 1;
      report "Test 3 FAILED TX. tx_sampled dec=" &
             integer'image(to_integer(unsigned(tx_sampled)))
        severity error;
    else
      report "Test 3 PASSED" severity note;
    end if;

    wait until falling_edge(sclk);
    wait for C_SCLK_PERIOD;  -- CS high ≥ 1 SCLK
    wait for C_SCLK_PERIOD;

    -------------------------------------------------------------------------
    -- Test 4: Multi-byte full-duplex, 3 bytes under one CS
    -------------------------------------------------------------------------
    report "Test 4: 3-byte full-duplex under single CS" severity note;

    -- prepare first TX byte, keep tx_valid high so PHY can sample at byte boundaries
    tx_valid <= '1';
    tx_byte  <= miso_seq(0);

    -- clear capture buffers
    for k in 0 to 3 loop
      mosi_captured(k) := (others => '0');
      miso_captured(k) := (others => '0');
    end loop;

    cs_n <= '0';
    -- 3 bytes, back-to-back, CS held low
    for j in 0 to 3 loop
      tx_byte <= miso_seq(j);
      spi_full_duplex(mosi_seq(j), miso_captured(j));
      -- Wait for rx_valid and settle
      wait until rx_valid = '1';
      --wait until falling_edge(sclk); 
      mosi_captured(j) := rx_byte;
    end loop;

    cs_n <= '1';
    tx_valid <= '0';
    wait for C_SCLK_PERIOD;  -- CS high ≥ 1 SCLK

    -- Check all three RX bytes
    for j in 0 to 3 loop
      if mosi_captured(j) /= mosi_seq(j) then
        error_count := error_count + 1;
        report "Test 4 FAILED RX byte " & integer'image(j) &
               " dec=" & integer'image(to_integer(unsigned(mosi_captured(j))))
          severity error;
      end if;
    end loop;

    -- Check all three TX bytes
    for j in 0 to 3 loop
      if miso_captured(j) /= miso_seq(j) then
        error_count := error_count + 1;
        report "Test 4 FAILED TX byte " & integer'image(j) &
               " dec=" & integer'image(to_integer(unsigned(miso_captured(j))))
          severity error;
      end if;
    end loop;

    if error_count = 0 then
      report "Test 4 PASSED" severity note;
    end if;


    -------------------------------------------------------------------------
    -- Summary
    -------------------------------------------------------------------------
    if error_count = 0 then
      report "All tests PASSED" severity note;
    else
      report "TESTBENCH FAILED, error_count=" &
             integer'image(error_count)
        severity error;
    end if;

    wait for 5*C_SCLK_PERIOD;
    wait;
  end process;

end architecture sim;
